# ====================================================================
#
#      usbs_eth.cdl
#
#      USB slave-side ethernet package.
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2003 Bart Veer
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      bartv
# Original data:  bartv
# Contributors:
# Date:           2000-10-04
#
#####DESCRIPTIONEND####
# ====================================================================

cdl_package CYGPKG_IO_USB_SLAVE_ETH {
    display     "USB slave ethernet support"
    include_dir "cyg/io/usb"
    parent      CYGPKG_IO_USB_SLAVE
    requires    { CYGHWR_IO_USB_SLAVE_OUT_ENDPOINTS >= 1 }
    requires    { CYGHWR_IO_USB_SLAVE_IN_ENDPOINTS >= 1 }
    compile     usbseth.c
    implements  CYGINT_IO_USB_SLAVE_CLIENTS
    doc         ref/io-usb-slave-eth.html
    
    description "
        The USB slave ethernet package supports the development
        of USB peripherals which provide an ethernet service to
        the host machine. Such a peripheral could be a simple
        USB-ethernet converter, or it could be rather more
        complicated internally."

    cdl_component CYGPKG_USBS_ETHDRV {
	display         "Provide a driver for a TCP/IP stack."
        requires        CYGPKG_IO_ETH_DRIVERS
	implements      CYGHWR_NET_DRIVERS
	default_value   CYGPKG_NET
	compile         -library=libextras.a usbsethdrv.c

	description "
	    The primary purpose of USB slave ethernet support is to provide
	    an ethernet service to the USB host. This is very different
	    from a conventional network driver which provides a service
            to a TCP/IP stack running inside the peripheral. If this
	    component is enabled then the USB-ethernet code will implement
	    an eCos network driver, thus supporting both a host-side TCP/IP
	    stack and an eCos stack. This raises issues such as enabling
	    the bridge code in the stack, and the package documentation
            should be consulted for further information."

	cdl_option CYGFUN_USBS_ETHDRV_STATISTICS {
	    display       "Maintain traffic statistics"
	    flavor        bool
	    default_value CYGPKG_SNMPAGENT
	    description "
	        The USB network device driver can maintain some statistics
                about traffic, for example the number of incoming and
	        outgoing packets. These statistics are intended mainly
	        for SNMP agent software."
	}

	cdl_option CYGDAT_USBS_ETHDRV_NAME {
	    display       "Name to use for this network device"
	    flavor        data
	    default_value { (1 == CYGHWR_NET_DRIVERS) ? "\"eth0\"" : "\"eth1\"" }
	    description "
	        The name of this network device for control purposes.
	    "
	}

	cdl_option CYGPRI_USBS_ETHDRV_ETH0 {
	    display       "Enable/disable generic eth0 configury"
	    flavor        bool
	    calculated    { "\"eth0\"" == CYGDAT_USBS_ETHDRV_NAME }
	    implements    CYGHWR_NET_DRIVER_ETH0
	    requires      !CYGHWR_NET_DRIVER_ETH0_BOOTP
	}
	
	cdl_option CYGPRI_USBS_ETHDRV_ETH1 {
	    display       "Enable/disable generic eth1 configury"
	    flavor        bool
	    calculated    { "\"eth1\"" == CYGDAT_USBS_ETHDRV_NAME }
	    implements    CYGHWR_NET_DRIVER_ETH1
	    requires      !CYGHWR_NET_DRIVER_ETH1_BOOTP
	}
    }
    
    cdl_component CYGPKG_IO_USB_SLAVE_ETH_OPTIONS {
	display     "Build options"
	flavor      none

	description "
	    Package-specific build options including control over compiler
	    flags used only in building this package."

	cdl_option CYGPKG_IO_USB_SLAVE_ETH_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building this package. These flags are used in addition
                to the set of global flags."
	}
        cdl_option CYGPKG_IO_USB_SLAVE_ETH_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building this package. These flags are removed from
                the set of global flags if present."
        }
    }
}
