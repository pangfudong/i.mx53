# ====================================================================
#
#      diagnosis.cdl
#
#      diagnosis configuration data. 
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2008 Freescale
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Fred.Fan
# Original data:  Fred.Fan
# Contributors:
# Date:           2008-03-15
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DIAGNOSIS {
    display       "Diagnostic tools"
    include_dir   cyg/diagnosis
#   doc           ref/services-diagnosis.html

    description "
      This package provides support for hardware diagnosis."

    compile -library=libextras.a core.c 

    cdl_component CYGPKG_MEMORY_DIAGNOSIS {
        display "memory diagnosis"
        flavor  bool

	description "This option includes memory test cases."
	
        compile -library=libextras.a memory/cmds.c
	
	cdl_option CYGSEM_RAM_RW_DIAGNOSIS {
                display "perform ram read/write diagnosis"
                flavor  bool
                default_value 1
         
	       	description      "
                    This option is overriden by the configuration in hal."

		compile memory/ram_rw.c
	}
    }
}


