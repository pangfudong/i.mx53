# ====================================================================
#
#      io_pci.cdl
#
#      eCos PCI library configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Contributors:
# Date:           1999-08-12
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_IO_PCI {
    display       "PCI configuration library"
    doc           ref/io-pci.html
    include_dir   cyg/io
    parent        CYGPKG_IO
    description   "
           The PCI configuration library provides initialization of devices
           on the PCI bus. Functions to find and access these devices are
	   also provided."

    compile       pci.c pci_hw.c

    cdl_component CYGPKG_IO_PCI_OPTIONS {
        display "PCI build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_IO_PCI_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the PCI configuration library. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_IO_PCI_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the PCI configuration library. These flags are removed from
                the set of global flags if present."
        }

        cdl_option CYGPKG_IO_PCI_DEBUG {
            display "Enable debugging."
            flavor  bool
            default_value 0
            description   "
                This option enables minimal debugging of the PCI library.
                In particular, it will print information about devices as the
                PCI bus is being scanned/searched."
        }

        cdl_option CYGPKG_IO_PCI_TESTS {
            display "PCI tests"
            flavor  data
            no_define
            calculated { "tests/pci1 tests/pci2" }
            description   "
                This option specifies the set of tests for the PCI configuration library."
        }

        cdl_option CYGPKG_IO_PCI_CONFIGURE_INTLINE {
            display "Writeback Interrupt Line register."
            flavor  bool
            default_value 0
            description   "
                This option causes a PCI device interrupt vector to be
                written to the Interrupt Line register in config space.
                This is traditionally done by a BIOS so that device
                drivers can read the interrupt vector directly from
                device configuration space."
        }
    }
}
