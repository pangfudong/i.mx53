# ====================================================================
#
#      ser_arm_aim711.cdl
#
#      eCos serial ARM Industrial Module AIM 711 configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Lars.Lindqvist@combitechsystems.com, rcassebohm
# Contributors:   jlarmour, rcassebohm
# Date:           2004-09-09
#
#####DESCRIPTIONEND####
#
# ====================================================================


cdl_package CYGPKG_IO_SERIAL_ARM_AIM711 {
    display       "ARM Industrial Module AIM 711 serial device drivers"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    active_if     CYGPKG_HAL_ARM_AIM711

    include_dir   cyg/io
    description   "
           This package contains serial device drivers for the
           ARM Industrial Module AIM 711."

    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#ifndef CYGDAT_IO_SERIAL_DEVICE_HEADER"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_DEVICE_HEADER <pkgconf/io_serial_arm_aim711.h>"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_GENERIC_16X5X_INL <cyg/io/ser_arm_aim711_16x5x.inl>"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_GENERIC_16X5X_CFG <pkgconf/io_serial_arm_aim711.h>"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_ARM_S3C4510_INL <cyg/io/ser_arm_aim711_s3c4510.inl>"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_ARM_S3C4510_CFG <pkgconf/io_serial_arm_aim711.h>"
        puts $::cdl_system_header "#endif"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
        puts $::cdl_header "#include <pkgconf/system.h>";
        puts $::cdl_header "#include <pkgconf/io_serial_arm_s3c4510.h>";
        puts $::cdl_header "#include <pkgconf/io_serial_generic_16x5x.h>";
    }

    cdl_component CYGPKG_IO_SERIAL_ARM_AIM711_16X5X {
        display       "ARM Industrial Module AIM 711 16x5x serial device drivers"

        parent        CYGPKG_IO_SERIAL_DEVICES
        active_if     CYGPKG_IO_SERIAL
        active_if     CYGPKG_HAL_ARM_AIM711
        default_value 1

        requires      CYGPKG_ERROR
        description   "
               This package contains serial device drivers for the
               ARM Industrial Module AIM 711 for the 16550 serial
               interface on board."

        # FIXME: This really belongs in the GENERIC_16X5X package
        cdl_interface CYGINT_IO_SERIAL_GENERIC_16X5X_REQUIRED {
            display   "Generic 16x5x serial driver required"
        }

        cdl_component CYGPKG_IO_SERIAL_ARM_AIM711_16X5X_SERIAL0 {
            display       "AIM 711 16X5X serial port 0 driver (COM1)"
            flavor        bool
            default_value 1
            description   "
                This option includes the serial device driver for the AIM 711 16X5X 
                port 0, which is COM1 on the AIM 711."

            implements    CYGINT_IO_SERIAL_GENERIC_16X5X_REQUIRED
            implements    CYGINT_IO_SERIAL_FLOW_CONTROL_HW
            implements    CYGINT_IO_SERIAL_LINE_STATUS_HW

            cdl_option CYGDAT_IO_SERIAL_ARM_AIM711_16X5X_SERIAL0_NAME {
                display       "Device name for the AIM 711 16X5X serial port 0 driver (COM1)"
                flavor        data
                default_value {"\"/dev/ser1\""}
                description   "
                    This option sets the name of the serial device for the AIM 711 
                    16X5X port 0 (COM1)."
            }

            cdl_option CYGNUM_IO_SERIAL_ARM_AIM711_16X5X_SERIAL0_BAUD {
                display       "Baud rate for the AIM 711 16X5X serial port 0 driver"
                flavor        data
                legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                              4800 7200 9600 14400 19200 38400 57600 115200 230400
                }
                default_value 38400
                description   "
                    This option specifies the default baud rate (speed) for the 
                    AIM 711 16X5X port 0."
            }

            cdl_option CYGNUM_IO_SERIAL_ARM_AIM711_16X5X_SERIAL0_BUFSIZE {
                display       "Buffer size for the AIM 711 16X5X serial port 0 driver"
                flavor        data
                legal_values  0 to 8192
                default_value 128
                description   "
                    This option specifies the size of the internal buffers used for
                    the AIM 711 16X5X port 0."
            }
        }
    }

    cdl_component CYGPKG_IO_SERIAL_ARM_AIM711_S3C4510 {
        display       "ARM Industrial Module AIM 711 S3C4510 serial device drivers"

        parent        CYGPKG_IO_SERIAL_DEVICES
        active_if     CYGPKG_IO_SERIAL
        active_if     CYGPKG_HAL_ARM_AIM711
        default_value 1

        requires      CYGPKG_ERROR
        description   "
               This package contains serial device drivers for the
               ARM Industrial Module AIM 711 for the internal serial
               interface of the S3C4510."

        # FIXME: This really belongs in the SERIAL_ARM_S3C4510 package
        cdl_interface CYGINT_IO_SERIAL_ARM_S3C4510_REQUIRED {
            display   "Generic s3c4510 serial driver required"
        }

        cdl_component CYGPKG_IO_SERIAL_ARM_AIM711_S3C4510_SERIAL0 {
            display       "AIM 711 S3C4510 serial port 0 driver (service adapter)"
            flavor        bool
            default_value 1
            description   "
                This option includes the serial device driver for the AIM 711 S3C4510 
                port 0, which is on the AIM 711 the port on the service adapter."

            implements    CYGINT_IO_SERIAL_ARM_S3C4510_REQUIRED

            cdl_option CYGDAT_IO_SERIAL_ARM_AIM711_S3C4510_SERIAL0_NAME {
                display       "Device name for the AIM 711 S3C4510 serial port 0 driver (service adapter)"
                flavor        data
                default_value {"\"/dev/ser0\""}
                description   "
                    This option sets the name of the serial device for the AIM 711 
                    S3C4510 port 0 (service adapter)."
            }

            cdl_option CYGNUM_IO_SERIAL_ARM_AIM711_S3C4510_SERIAL0_BAUD {
                display       "Baud rate for the AIM 711 S3C4510 serial port 0 driver"
                flavor        data
                legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                              4800 7200 9600 14400 19200 38400 57600 115200 230400
                }
                default_value 38400
                description   "
                    This option specifies the default baud rate (speed) for the 
                    AIM 711 S3C4510 port 0."
            }

            cdl_option CYGNUM_IO_SERIAL_ARM_AIM711_S3C4510_SERIAL0_BUFSIZE {
                display       "Buffer size for the AIM 711 S3C4510 serial port 0 driver"
                flavor        data
                legal_values  0 to 8192
                default_value 128
                description   "
                    This option specifies the size of the internal buffers used for
                    the AIM 711 S3C4510 port 0."
            }
        }

        cdl_component CYGPKG_IO_SERIAL_ARM_AIM711_S3C4510_SERIAL1 {
            display       "AIM 711 S3C4510 serial port 1 driver (COM2)"
            flavor        bool
            default_value 1
            description   "
                This option includes the serial device driver for the AIM 711 
                S3C4510 port 1, which is the COM2 on the AIM 711."

            implements    CYGINT_IO_SERIAL_ARM_S3C4510_REQUIRED

            cdl_option CYGDAT_IO_SERIAL_ARM_AIM711_S3C4510_SERIAL1_NAME {
                display       "Device name for the AIM 711 S3C4510 serial port 1 driver (COM2)"
                flavor        data
                default_value {"\"/dev/ser2\""}
                description   "
                    This option specifies the name of serial device for the 
                    AIM 711 S3C4510 port 1 (COM2)."
            }

            cdl_option CYGNUM_IO_SERIAL_ARM_AIM711_S3C4510_SERIAL1_BAUD {
                display       "Baud rate for the AIM 711 S3C4510 serial port 1 driver"
                flavor        data
                legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                              4800 7200 9600 14400 19200 38400 57600 115200 230400
                }
                default_value 38400
                description   "
                    This option specifies the default baud rate (speed) for the 
                    AIM 711 S3C4510 port 1."
            }

            cdl_option CYGNUM_IO_SERIAL_ARM_AIM711_S3C4510_SERIAL1_BUFSIZE {
                display       "Buffer size for the AIM 711 S3C4510 serial port 1 driver"
                flavor        data
                legal_values  0 to 8192
                default_value 128
                description   "
                    This option specifies the size of the internal buffers used 
                    for the AIM 711 S3C4510 port 1."
            }
        }
    }

    cdl_component CYGPKG_IO_SERIAL_ARM_AIM711_OPTIONS {
        display "Serial device driver build options"
        flavor  none
        description   "
        Package specific build options including control over
        compiler flags used only in building this package,
        and details of which tests are built."


        cdl_option CYGPKG_IO_SERIAL_ARM_AIM711_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_IO_SERIAL_ARM_AIM711_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are removed from
                the set of global flags if present."
        }
    }

    cdl_component CYGPKG_IO_SERIAL_ARM_AIM711_TESTING {
        display    "Testing parameters"
        flavor     bool
        calculated 1
        active_if  CYGPKG_IO_SERIAL_ARM_AIM711_16X5X_SERIAL0

        cdl_option CYGPRI_SER_TEST_SER_DEV {
            display       "Serial device used for testing"
            flavor        data
            default_value { CYGDAT_IO_SERIAL_ARM_AIM711_16X5X_SERIAL0_NAME }
        }

        define_proc {
            puts $::cdl_header "#define CYGPRI_SER_TEST_CRASH_ID \"arm16x5x\""
            puts $::cdl_header "#define CYGPRI_SER_TEST_TTY_DEV  \"/dev/tty2\""
        }
    }
}

# EOF ser_arm_aim711.cdl
