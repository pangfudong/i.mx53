# ====================================================================
#
#      blib.cdl
#
#      Block cache and access library configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2003 Savin Zlobec 
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      savin 
# Contributors:   
# Date:           2003-08-29
#
#####DESCRIPTIONEND####
# ====================================================================

cdl_package CYGPKG_BLOCK_LIB {
    display         "Block cache and access library"
    define_header   blib.h
    include_dir     blib

    requires        CYGPKG_ISOINFRA
    requires        CYGPKG_MEMALLOC
    requires        CYGPKG_LINUX_COMPAT
    requires        CYGPKG_ERROR
    
    compile         -library=libextras.a blib.c    

    cdl_option CYGIMP_BLOCK_LIB_STATISTICS {
        display         "Block access statistics support"
        flavor          bool
        default_value   1
        description     "This option enables statistics for
                         block access operations."
    }
}

# ====================================================================
# End of blib.cdl
