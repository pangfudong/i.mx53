# ====================================================================
#
#      ide_disk.cdl
#
#      A generic IDE disk driver package.
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2004 Red Hat, Inc.
## Copyright (C) 2004 eCosCentric, Ltd
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      iz
# Contributors:
# Date:           2004-10-16
#
#####DESCRIPTIONEND####
# ====================================================================

cdl_package CYGPKG_DEVS_DISK_IDE {
    display     "Disk driver for generic IDE"
    
    parent      CYGPKG_IO_DISK_DEVICES
    active_if   CYGPKG_IO_DISK

    compile     -library=libextras.a   ide_disk.c
    
    cdl_component CYGVAR_DEVS_DISK_IDE_DISK0 {
    	display         "Provide disk 0 device"
        flavor          bool
        default_value   1
        description     "IDE chanel 0:0 disk driver"
        
        cdl_option CYGDAT_IO_DISK_IDE_DISK0_NAME {
            display       "Device name for disk 0 device"
            flavor        data
            default_value {"\"/dev/hda/\""}
        }
    }
    
    cdl_component CYGVAR_DEVS_DISK_IDE_DISK1 {
     display         "Provide disk 1 device"
        flavor          bool
        default_value   0
        description     "IDE chanel 0:1 disk driver"
        
        cdl_option CYGDAT_IO_DISK_IDE_DISK1_NAME {
            display       "Device name for disk 1 device"
            flavor        data
            default_value {"\"/dev/hdb/\""}
        }
    }
    
    cdl_component CYGVAR_DEVS_DISK_IDE_DISK2 {
     display         "Provide disk 2 device"
        flavor          bool
        default_value   0
        description     "IDE chanel 1:0 disk driver"
        
        cdl_option CYGDAT_IO_DISK_IDE_DISK2_NAME {
            display       "Device name for disk 2 device"
            flavor        data
            default_value {"\"/dev/hdc/\""}
        }
    }
    
    cdl_component CYGVAR_DEVS_DISK_IDE_DISK3 {
     display         "Provide disk 3 device"
        flavor          bool
        default_value   0
        description     "IDE chanel 1:1 disk driver"
        
        cdl_option CYGDAT_IO_DISK_IDE_DISK3_NAME {
            display       "Device name for disk 3 device"
            flavor        data
            default_value {"\"/dev/hdd/\""}
        }
    }

    cdl_option CYGDAT_DEVS_DISK_IDE_SECTOR_SIZE {
        display       "Disk sector size"
        flavor        data
        default_value 512
        description "
        This option controls the disk sector size (default=512)"
     }

    cdl_option CYGSEM_DEVS_DISK_IDE_VMWARE {
        display       "Work with VMware virtual disks"
        flavor        bool
        default_value 0
        description "
        This option controls the disk driver behaviour at ide-init"
     }

}

# EOF ide_disk.cdl
