# ====================================================================
#
#      flash_toshiba_tc58xxx.cdl
#
#      FLASH memory - Hardware support for Toshiba TC58xxx parts
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
## Copyright (C) 2003 Gary Thomas
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Gary Thomas <gary@mlbassoc.com>
# Contributors:   
# Date:           2003-09-02
# Description:    FLASH drivers for Toshiba TC58xxx NAND devices.  Based on
#                 Atmel AT49xxxx drivers by Jani Monoses <jani@iv.ro>
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_TOSHIBA_TC58XXX {
    display       "Toshiba TC58XXX FLASH memory support"
    description   "FLASH memory device support for Toshiba TC58XXX"
    parent        CYGPKG_IO_FLASH
    active_if	  CYGPKG_IO_FLASH
    requires      { CYGSEM_IO_FLASH_READ_INDIRECT == 1 }

    active_if     CYGINT_DEVS_FLASH_TOSHIBA_TC58XXX_REQUIRED

    implements    CYGHWR_IO_FLASH_DEVICE

    include_dir   cyg/io
}

# EOF flash_toshiba_tc58xxx.cdl
