# ====================================================================
#
#      sntp.cdl
#
#      Simple Network Time Protocol
#
# ====================================================================
######ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2003 Andrew Lunn
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
######ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Andrew Lunn
# Contributors:
# Date:           2003-02-11
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_NET_SNTP {
    display       "Simple Network Time Protocol Client (SNTP)"
    description   "
           This package provides a SNTP client which can recieve broadcast time 
           information and set the system clock."
    doc           ref/net-sntp.html
    include_dir   cyg/sntp

    requires      CYGPKG_NET
    requires      CYGPKG_LIBC_TIME
    requires      CYGSEM_LIBC_TIME_TIME_WORKING
    requires      CYGSEM_LIBC_TIME_SETTIME_WORKING
    compile       sntp.c
    
    cdl_component CYGPKG_NET_SNTP_UNICAST {
        display "Enable SNTP client unicast support"
        flavor  bool
        default_value 0
        description   "
            This option enables SNTP unicast mode in
            for the SNTP client.  This mode will send
            SNTP requests to NTP/SNTP servers in
            addition to listening for SNTP broadcasts."

        cdl_option CYGNUM_NET_SNTP_UNICAST_MAXDHCP {
            display "Maximum number of NTP servers to use from DHCP"
            flavor  booldata
            requires CYGPKG_NET_DHCP
            legal_values 1 to 8
            default_value 2
            description   "
                This option specifies the maximum number of
                NTP servers to get from DHCP.  These servers
                are used to configure the unicast SNTP client.
                Disabling this option disables DHCP usage."
        }
    }

    cdl_component CYGPKG_NET_SNTP_OPTIONS {
        display "SNTP support build options"
        flavor  none
        no_define

        cdl_option CYGPKG_NET_SNTP_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the SNTP package.
                These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_NET_SNTP_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the SNTP package. These flags are removed from
                the set of global flags if present."
        }
    }

    cdl_option CYGPKG_NET_SNTP_TESTS {
        display "sntp tests"
        flavor  data
        no_define
        calculated { CYGPKG_NET_BUILD_HW_TESTS ? "tests/sntp1.c" : "" }
    }
}

# ====================================================================
# EOF sntp.cdl
