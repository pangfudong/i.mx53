# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Original data:  gthomas
# Contributors:
# Date:           2000-07-26
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_ONMXC {
    display       "Support FLASH memory on Freescale MXC platforms"

    implements    CYGHWR_IO_FLASH_DEVICE
    parent        CYGPKG_IO_FLASH
    active_if	  CYGPKG_IO_FLASH

    include_dir   cyg/io

    cdl_option CYGHWR_DEVS_FLASH_MXC_NOR {
        display       "MXC platform NOR flash memory support"
        default_value 0
        description   "
            When this option is enabled, it indicates NOR flash is 
            supported on the MXC platforms"
        define_proc {
            puts $::cdl_system_header "#define MXCFLASH_SELECT_NOR"
        }
    }
    cdl_option CYGHWR_DEVS_FLASH_MXC_NAND {
        display       "MXC platform NAND flash memory support"
        default_value 0
        requires      { CYGSEM_IO_FLASH_READ_INDIRECT == 1 }
        description   "
            When this option is enabled, it indicates NAND flash is 
            supported on the MXC platforms"
        define_proc {
            puts $::cdl_system_header "#define MXCFLASH_SELECT_NAND"
        }
        compile       mxc_nfc.c
    }
    cdl_option CYGHWR_DEVS_FLASH_MXC_MULTI {
        display       "MXC platform multi flash memory support"
        default_value 1
        active_if     {CYGHWR_DEVS_FLASH_MXC_NAND && CYGHWR_DEVS_FLASH_MXC_NOR}
        description   "
            When this option is enabled, it indicates multi flashes are 
            supported on the MXC platforms (like NAND and NOR)"
        define_proc {
            puts $::cdl_system_header "#define MXCFLASH_SELECT_MULTI"
        }
        compile       mxcflash_wrapper.c
    }
    cdl_interface CYGHWR_DEVS_FLASH_MXC_NAND_RESET_WORKAROUND {
        display       "MXC platform NAND flash reset workaround support"
        active_if     {CYGHWR_DEVS_FLASH_MXC_NAND}
        description   "
            When this option is enabled, it indicates 0xFFFF is used for
            the NAND reset command instead of 0xFF."
    }
}